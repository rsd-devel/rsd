

localparam LED_WIDTH = 8;

`include "XilinxMacros.vh"

module RSD(
input
    wire clk,
    wire negResetIn,
output
    wire [LED_WIDTH-1:0] ledOut,
input
    wire  axi4MemoryIF_M_AXI_ACLK,
    wire  axi4MemoryIF_M_AXI_ARESETN,
output
    wire [1 : 0] axi4MemoryIF_M_AXI_AWID,
    wire [31 : 0] axi4MemoryIF_M_AXI_AWADDR,
    wire [7 : 0] axi4MemoryIF_M_AXI_AWLEN,
    wire [2 : 0] axi4MemoryIF_M_AXI_AWSIZE,
    wire [1 : 0] axi4MemoryIF_M_AXI_AWBURST,
    wire  axi4MemoryIF_M_AXI_AWLOCK,
    wire [3 : 0] axi4MemoryIF_M_AXI_AWCACHE,
    wire [2 : 0] axi4MemoryIF_M_AXI_AWPROT,
    wire [3 : 0] axi4MemoryIF_M_AXI_AWQOS,
    wire [0 : 1] axi4MemoryIF_M_AXI_AWUSER,
    wire  axi4MemoryIF_M_AXI_AWVALID,
input
    wire  axi4MemoryIF_M_AXI_AWREADY,
output
    wire [63 : 0] axi4MemoryIF_M_AXI_WDATA,
    wire [7 : 0] axi4MemoryIF_M_AXI_WSTRB,
    wire  axi4MemoryIF_M_AXI_WLAST,
    wire [0 : 1] axi4MemoryIF_M_AXI_WUSER,
    wire  axi4MemoryIF_M_AXI_WVALID,
input
    wire  axi4MemoryIF_M_AXI_WREADY,
    wire [1 : 0] axi4MemoryIF_M_AXI_BID,
    wire [1 : 0] axi4MemoryIF_M_AXI_BRESP,
    wire [0 : 1] axi4MemoryIF_M_AXI_BUSER,
    wire  axi4MemoryIF_M_AXI_BVALID,
output
    wire  axi4MemoryIF_M_AXI_BREADY,
    wire [1 : 0] axi4MemoryIF_M_AXI_ARID,
    wire [31 : 0] axi4MemoryIF_M_AXI_ARADDR,
    wire [7 : 0] axi4MemoryIF_M_AXI_ARLEN,
    wire [2 : 0] axi4MemoryIF_M_AXI_ARSIZE,
    wire [1 : 0] axi4MemoryIF_M_AXI_ARBURST,
    wire  axi4MemoryIF_M_AXI_ARLOCK,
    wire [3 : 0] axi4MemoryIF_M_AXI_ARCACHE,
    wire [2 : 0] axi4MemoryIF_M_AXI_ARPROT,
    wire [3 : 0] axi4MemoryIF_M_AXI_ARQOS,
    wire [0 : 1] axi4MemoryIF_M_AXI_ARUSER,
    wire  axi4MemoryIF_M_AXI_ARVALID,
input
    wire  axi4MemoryIF_M_AXI_ARREADY,
    wire [1 : 0] axi4MemoryIF_M_AXI_RID,
    wire [63 : 0] axi4MemoryIF_M_AXI_RDATA,
    wire [1 : 0] axi4MemoryIF_M_AXI_RRESP,
    wire  axi4MemoryIF_M_AXI_RLAST,
    wire [0 : 1] axi4MemoryIF_M_AXI_RUSER,
    wire  axi4MemoryIF_M_AXI_RVALID,
output
    wire  axi4MemoryIF_M_AXI_RREADY,
input
    wire axi4LitePlToPsControlRegisterIF_S_AXI_ACLK,
    wire axi4LitePlToPsControlRegisterIF_S_AXI_ARESETN,
    wire [6 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_ARADDR,
    wire [2 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_ARPROT,
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_ARVALID,
output
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_ARREADY,
    wire [31 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_RDATA,
    wire [1 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_RRESP,
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_RVALID,
input
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_RREADY,
    wire axi4LitePsToPlControlRegisterIF_S_AXI_ACLK,
    wire axi4LitePsToPlControlRegisterIF_S_AXI_ARESETN,
    wire [6 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_AWADDR,
    wire [2 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_AWPROT,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_AWVALID,
output
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_AWREADY,
input
    wire [31 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_WDATA,
    wire [3 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_WSTRB,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_WVALID,
output
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_WREADY,
    wire [1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_BRESP,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_BVALID,
input
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_BREADY,
    wire [6 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_ARADDR,
    wire [2 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_ARPROT,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_ARVALID,
output
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_ARREADY,
    wire [31 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_RDATA,
    wire [1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_RRESP,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_RVALID,
input
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_RREADY
);

    Main_Zynq_Wrapper main(
        .clk (clk),
        .negResetIn (negResetIn),
        .ledOut (ledOut),
        .axi4MemoryIF_M_AXI_ACLK (axi4MemoryIF_M_AXI_ACLK),
        .axi4MemoryIF_M_AXI_ARESETN (axi4MemoryIF_M_AXI_ARESETN),
        .axi4MemoryIF_M_AXI_AWID (axi4MemoryIF_M_AXI_AWID),
        .axi4MemoryIF_M_AXI_AWADDR (axi4MemoryIF_M_AXI_AWADDR),
        .axi4MemoryIF_M_AXI_AWLEN (axi4MemoryIF_M_AXI_AWLEN),
        .axi4MemoryIF_M_AXI_AWSIZE (axi4MemoryIF_M_AXI_AWSIZE),
        .axi4MemoryIF_M_AXI_AWBURST (axi4MemoryIF_M_AXI_AWBURST),
        .axi4MemoryIF_M_AXI_AWLOCK (axi4MemoryIF_M_AXI_AWLOCK),
        .axi4MemoryIF_M_AXI_AWCACHE (axi4MemoryIF_M_AXI_AWCACHE),
        .axi4MemoryIF_M_AXI_AWPROT (axi4MemoryIF_M_AXI_AWPROT),
        .axi4MemoryIF_M_AXI_AWQOS (axi4MemoryIF_M_AXI_AWQOS),
        .axi4MemoryIF_M_AXI_AWUSER (axi4MemoryIF_M_AXI_AWUSER),
        .axi4MemoryIF_M_AXI_AWVALID (axi4MemoryIF_M_AXI_AWVALID),
        .axi4MemoryIF_M_AXI_AWREADY (axi4MemoryIF_M_AXI_AWREADY),
        .axi4MemoryIF_M_AXI_WDATA (axi4MemoryIF_M_AXI_WDATA),
        .axi4MemoryIF_M_AXI_WSTRB (axi4MemoryIF_M_AXI_WSTRB),
        .axi4MemoryIF_M_AXI_WLAST (axi4MemoryIF_M_AXI_WLAST),
        .axi4MemoryIF_M_AXI_WUSER (axi4MemoryIF_M_AXI_WUSER),
        .axi4MemoryIF_M_AXI_WVALID (axi4MemoryIF_M_AXI_WVALID),
        .axi4MemoryIF_M_AXI_WREADY (axi4MemoryIF_M_AXI_WREADY),
        .axi4MemoryIF_M_AXI_BID (axi4MemoryIF_M_AXI_BID),
        .axi4MemoryIF_M_AXI_BRESP (axi4MemoryIF_M_AXI_BRESP),
        .axi4MemoryIF_M_AXI_BUSER (axi4MemoryIF_M_AXI_BUSER),
        .axi4MemoryIF_M_AXI_BVALID (axi4MemoryIF_M_AXI_BVALID),
        .axi4MemoryIF_M_AXI_BREADY (axi4MemoryIF_M_AXI_BREADY),
        .axi4MemoryIF_M_AXI_ARID (axi4MemoryIF_M_AXI_ARID),
        .axi4MemoryIF_M_AXI_ARADDR (axi4MemoryIF_M_AXI_ARADDR),
        .axi4MemoryIF_M_AXI_ARLEN (axi4MemoryIF_M_AXI_ARLEN),
        .axi4MemoryIF_M_AXI_ARSIZE (axi4MemoryIF_M_AXI_ARSIZE),
        .axi4MemoryIF_M_AXI_ARBURST (axi4MemoryIF_M_AXI_ARBURST),
        .axi4MemoryIF_M_AXI_ARLOCK (axi4MemoryIF_M_AXI_ARLOCK),
        .axi4MemoryIF_M_AXI_ARCACHE (axi4MemoryIF_M_AXI_ARCACHE),
        .axi4MemoryIF_M_AXI_ARPROT (axi4MemoryIF_M_AXI_ARPROT),
        .axi4MemoryIF_M_AXI_ARQOS (axi4MemoryIF_M_AXI_ARQOS),
        .axi4MemoryIF_M_AXI_ARUSER (axi4MemoryIF_M_AXI_ARUSER),
        .axi4MemoryIF_M_AXI_ARVALID (axi4MemoryIF_M_AXI_ARVALID),
        .axi4MemoryIF_M_AXI_ARREADY (axi4MemoryIF_M_AXI_ARREADY),
        .axi4MemoryIF_M_AXI_RID (axi4MemoryIF_M_AXI_RID),
        .axi4MemoryIF_M_AXI_RDATA (axi4MemoryIF_M_AXI_RDATA),
        .axi4MemoryIF_M_AXI_RRESP (axi4MemoryIF_M_AXI_RRESP),
        .axi4MemoryIF_M_AXI_RLAST (axi4MemoryIF_M_AXI_RLAST),
        .axi4MemoryIF_M_AXI_RUSER (axi4MemoryIF_M_AXI_RUSER),
        .axi4MemoryIF_M_AXI_RVALID (axi4MemoryIF_M_AXI_RVALID),
        .axi4MemoryIF_M_AXI_RREADY (axi4MemoryIF_M_AXI_RREADY),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ACLK (axi4LitePlToPsControlRegisterIF_S_AXI_ACLK),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARESETN (axi4LitePlToPsControlRegisterIF_S_AXI_ARESETN),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARADDR (axi4LitePlToPsControlRegisterIF_S_AXI_ARADDR),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARPROT (axi4LitePlToPsControlRegisterIF_S_AXI_ARPROT),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARVALID (axi4LitePlToPsControlRegisterIF_S_AXI_ARVALID),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARREADY (axi4LitePlToPsControlRegisterIF_S_AXI_ARREADY),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RDATA (axi4LitePlToPsControlRegisterIF_S_AXI_RDATA),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RRESP (axi4LitePlToPsControlRegisterIF_S_AXI_RRESP),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RVALID (axi4LitePlToPsControlRegisterIF_S_AXI_RVALID),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RREADY (axi4LitePlToPsControlRegisterIF_S_AXI_RREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ACLK (axi4LitePsToPlControlRegisterIF_S_AXI_ACLK),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARESETN (axi4LitePsToPlControlRegisterIF_S_AXI_ARESETN),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWADDR (axi4LitePsToPlControlRegisterIF_S_AXI_AWADDR),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWPROT (axi4LitePsToPlControlRegisterIF_S_AXI_AWPROT),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWVALID (axi4LitePsToPlControlRegisterIF_S_AXI_AWVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWREADY (axi4LitePsToPlControlRegisterIF_S_AXI_AWREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WDATA (axi4LitePsToPlControlRegisterIF_S_AXI_WDATA),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WSTRB (axi4LitePsToPlControlRegisterIF_S_AXI_WSTRB),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WVALID (axi4LitePsToPlControlRegisterIF_S_AXI_WVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WREADY (axi4LitePsToPlControlRegisterIF_S_AXI_WREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_BRESP (axi4LitePsToPlControlRegisterIF_S_AXI_BRESP),
        .axi4LitePsToPlControlRegisterIF_S_AXI_BVALID (axi4LitePsToPlControlRegisterIF_S_AXI_BVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_BREADY (axi4LitePsToPlControlRegisterIF_S_AXI_BREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARADDR (axi4LitePsToPlControlRegisterIF_S_AXI_ARADDR),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARPROT (axi4LitePsToPlControlRegisterIF_S_AXI_ARPROT),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARVALID (axi4LitePsToPlControlRegisterIF_S_AXI_ARVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARREADY (axi4LitePsToPlControlRegisterIF_S_AXI_ARREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RDATA (axi4LitePsToPlControlRegisterIF_S_AXI_RDATA),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RRESP (axi4LitePsToPlControlRegisterIF_S_AXI_RRESP),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RVALID (axi4LitePsToPlControlRegisterIF_S_AXI_RVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RREADY (axi4LitePsToPlControlRegisterIF_S_AXI_RREADY)
    );

endmodule : RSD
