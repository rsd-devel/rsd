
`include "SysDeps/XilinxMacros.vh"

localparam LED_WIDTH = 8;

module RSD(
input
    wire clk,
    wire negResetIn,
output
    wire [LED_WIDTH-1:0] ledOut,
input
    wire  axi4MemoryIF_M_AXI_ACLK,
    wire  axi4MemoryIF_M_AXI_ARESETN,
output
    wire [`MEMORY_AXI4_WRITE_ID_WIDTH-1 : 0] axi4MemoryIF_M_AXI_AWID,
    wire [`MEMORY_AXI4_ADDR_BIT_SIZE-1 : 0] axi4MemoryIF_M_AXI_AWADDR,
    wire [`MEMORY_AXI4_AWLEN_WIDTH-1 : 0] axi4MemoryIF_M_AXI_AWLEN,
    wire [`MEMORY_AXI4_AWSIZE_WIDTH-1 : 0] axi4MemoryIF_M_AXI_AWSIZE,
    wire [`MEMORY_AXI4_AWBURST_WIDTH-1 : 0] axi4MemoryIF_M_AXI_AWBURST,
    wire  axi4MemoryIF_M_AXI_AWLOCK,
    wire [`MEMORY_AXI4_AWCACHE_WIDTH-1 : 0] axi4MemoryIF_M_AXI_AWCACHE,
    wire [`MEMORY_AXI4_AWPROT_WIDTH-1 : 0] axi4MemoryIF_M_AXI_AWPROT,
    wire [`MEMORY_AXI4_AWQOS_WIDTH-1 : 0] axi4MemoryIF_M_AXI_AWQOS,
    wire [`MEMORY_AXI4_AWUSER_WIDTH-1 : 1] axi4MemoryIF_M_AXI_AWUSER,
    wire  axi4MemoryIF_M_AXI_AWVALID,
input
    wire  axi4MemoryIF_M_AXI_AWREADY,
output
    wire [`MEMORY_AXI4_DATA_BIT_NUM-1 : 0] axi4MemoryIF_M_AXI_WDATA,
    wire [`MEMORY_AXI4_DATA_BIT_NUM/8-1 : 0] axi4MemoryIF_M_AXI_WSTRB,
    wire  axi4MemoryIF_M_AXI_WLAST,
    wire [`MEMORY_AXI4_WUSER_WIDTH-1 : 1] axi4MemoryIF_M_AXI_WUSER,
    wire  axi4MemoryIF_M_AXI_WVALID,
input
    wire  axi4MemoryIF_M_AXI_WREADY,
    wire [`MEMORY_AXI4_WRITE_ID_WIDTH-1 : 0] axi4MemoryIF_M_AXI_BID,
    wire [`MEMORY_AXI4_BRESP_WIDTH-1 : 0] axi4MemoryIF_M_AXI_BRESP,
    wire [`MEMORY_AXI4_BUSER_WIDTH-1 : 0] axi4MemoryIF_M_AXI_BUSER,
    wire  axi4MemoryIF_M_AXI_BVALID,
output
    wire  axi4MemoryIF_M_AXI_BREADY,
    wire [`MEMORY_AXI4_READ_ID_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARID,
    wire [`MEMORY_AXI4_ADDR_BIT_SIZE-1 : 0] axi4MemoryIF_M_AXI_ARADDR,
    wire [`MEMORY_AXI4_ARLEN_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARLEN,
    wire [`MEMORY_AXI4_ARSIZE_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARSIZE,
    wire [`MEMORY_AXI4_ARBURST_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARBURST,
    wire  axi4MemoryIF_M_AXI_ARLOCK,
    wire [`MEMORY_AXI4_ARCACHE_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARCACHE,
    wire [`MEMORY_AXI4_ARPROT_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARPROT,
    wire [`MEMORY_AXI4_ARQOS_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARQOS,
    wire [`MEMORY_AXI4_ARUSER_WIDTH-1 : 0] axi4MemoryIF_M_AXI_ARUSER,
    wire  axi4MemoryIF_M_AXI_ARVALID,
input
    wire  axi4MemoryIF_M_AXI_ARREADY,
    wire [`MEMORY_AXI4_READ_ID_WIDTH-1 : 0] axi4MemoryIF_M_AXI_RID,
    wire [`MEMORY_AXI4_DATA_BIT_NUM-1 : 0] axi4MemoryIF_M_AXI_RDATA,
    wire [`MEMORY_AXI4_RRESP_WIDTH-1 : 0] axi4MemoryIF_M_AXI_RRESP,
    wire  axi4MemoryIF_M_AXI_RLAST,
    wire [`MEMORY_AXI4_RUSER_WIDTH-1 : 0] axi4MemoryIF_M_AXI_RUSER,
    wire  axi4MemoryIF_M_AXI_RVALID,
output
    wire  axi4MemoryIF_M_AXI_RREADY,
input
    wire axi4LitePlToPsControlRegisterIF_S_AXI_ACLK,
    wire axi4LitePlToPsControlRegisterIF_S_AXI_ARESETN,
    wire [`PS_PL_CTRL_REG_ADDR_BIT_SIZE-1 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_ARADDR,
    wire [`PS_PL_CTRL_REG_AWPROT_WIDTH-1 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_ARPROT,
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_ARVALID,
output
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_ARREADY,
    wire [`PS_PL_CTRL_REG_DATA_BIT_SIZE-1 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_RDATA,
    wire [`PS_PL_CTRL_REG_RRESP_WIDTH-1 : 0] axi4LitePlToPsControlRegisterIF_S_AXI_RRESP,
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_RVALID,
input
    wire  axi4LitePlToPsControlRegisterIF_S_AXI_RREADY,
    wire axi4LitePsToPlControlRegisterIF_S_AXI_ACLK,
    wire axi4LitePsToPlControlRegisterIF_S_AXI_ARESETN,
    wire [`PS_PL_CTRL_REG_ADDR_BIT_SIZE-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_AWADDR,
    wire [`PS_PL_CTRL_REG_AWPROT_WIDTH-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_AWPROT,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_AWVALID,
output
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_AWREADY,
input
    wire [`PS_PL_CTRL_REG_DATA_BIT_SIZE-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_WDATA,
    wire [(`PS_PL_CTRL_REG_DATA_BIT_SIZE/8)-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_WSTRB,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_WVALID,
output
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_WREADY,
    wire [`PS_PL_CTRL_REG_BRESP_WIDTH-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_BRESP,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_BVALID,
input
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_BREADY,
    wire [`PS_PL_CTRL_REG_ADDR_BIT_SIZE-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_ARADDR,
    wire [`PS_PL_CTRL_REG_ARPROT_WIDTH-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_ARPROT,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_ARVALID,
output
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_ARREADY,
    wire [`PS_PL_CTRL_REG_DATA_BIT_SIZE-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_RDATA,
    wire [`PS_PL_CTRL_REG_RRESP_WIDTH-1 : 0] axi4LitePsToPlControlRegisterIF_S_AXI_RRESP,
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_RVALID,
input
    wire  axi4LitePsToPlControlRegisterIF_S_AXI_RREADY
);

    Main_Zynq_Wrapper main(
        .clk (clk),
        .negResetIn (negResetIn),
        .ledOut (ledOut),
        .axi4MemoryIF_M_AXI_ACLK (axi4MemoryIF_M_AXI_ACLK),
        .axi4MemoryIF_M_AXI_ARESETN (axi4MemoryIF_M_AXI_ARESETN),
        .axi4MemoryIF_M_AXI_AWID (axi4MemoryIF_M_AXI_AWID),
        .axi4MemoryIF_M_AXI_AWADDR (axi4MemoryIF_M_AXI_AWADDR),
        .axi4MemoryIF_M_AXI_AWLEN (axi4MemoryIF_M_AXI_AWLEN),
        .axi4MemoryIF_M_AXI_AWSIZE (axi4MemoryIF_M_AXI_AWSIZE),
        .axi4MemoryIF_M_AXI_AWBURST (axi4MemoryIF_M_AXI_AWBURST),
        .axi4MemoryIF_M_AXI_AWLOCK (axi4MemoryIF_M_AXI_AWLOCK),
        .axi4MemoryIF_M_AXI_AWCACHE (axi4MemoryIF_M_AXI_AWCACHE),
        .axi4MemoryIF_M_AXI_AWPROT (axi4MemoryIF_M_AXI_AWPROT),
        .axi4MemoryIF_M_AXI_AWQOS (axi4MemoryIF_M_AXI_AWQOS),
        .axi4MemoryIF_M_AXI_AWUSER (axi4MemoryIF_M_AXI_AWUSER),
        .axi4MemoryIF_M_AXI_AWVALID (axi4MemoryIF_M_AXI_AWVALID),
        .axi4MemoryIF_M_AXI_AWREADY (axi4MemoryIF_M_AXI_AWREADY),
        .axi4MemoryIF_M_AXI_WDATA (axi4MemoryIF_M_AXI_WDATA),
        .axi4MemoryIF_M_AXI_WSTRB (axi4MemoryIF_M_AXI_WSTRB),
        .axi4MemoryIF_M_AXI_WLAST (axi4MemoryIF_M_AXI_WLAST),
        .axi4MemoryIF_M_AXI_WUSER (axi4MemoryIF_M_AXI_WUSER),
        .axi4MemoryIF_M_AXI_WVALID (axi4MemoryIF_M_AXI_WVALID),
        .axi4MemoryIF_M_AXI_WREADY (axi4MemoryIF_M_AXI_WREADY),
        .axi4MemoryIF_M_AXI_BID (axi4MemoryIF_M_AXI_BID),
        .axi4MemoryIF_M_AXI_BRESP (axi4MemoryIF_M_AXI_BRESP),
        .axi4MemoryIF_M_AXI_BUSER (axi4MemoryIF_M_AXI_BUSER),
        .axi4MemoryIF_M_AXI_BVALID (axi4MemoryIF_M_AXI_BVALID),
        .axi4MemoryIF_M_AXI_BREADY (axi4MemoryIF_M_AXI_BREADY),
        .axi4MemoryIF_M_AXI_ARID (axi4MemoryIF_M_AXI_ARID),
        .axi4MemoryIF_M_AXI_ARADDR (axi4MemoryIF_M_AXI_ARADDR),
        .axi4MemoryIF_M_AXI_ARLEN (axi4MemoryIF_M_AXI_ARLEN),
        .axi4MemoryIF_M_AXI_ARSIZE (axi4MemoryIF_M_AXI_ARSIZE),
        .axi4MemoryIF_M_AXI_ARBURST (axi4MemoryIF_M_AXI_ARBURST),
        .axi4MemoryIF_M_AXI_ARLOCK (axi4MemoryIF_M_AXI_ARLOCK),
        .axi4MemoryIF_M_AXI_ARCACHE (axi4MemoryIF_M_AXI_ARCACHE),
        .axi4MemoryIF_M_AXI_ARPROT (axi4MemoryIF_M_AXI_ARPROT),
        .axi4MemoryIF_M_AXI_ARQOS (axi4MemoryIF_M_AXI_ARQOS),
        .axi4MemoryIF_M_AXI_ARUSER (axi4MemoryIF_M_AXI_ARUSER),
        .axi4MemoryIF_M_AXI_ARVALID (axi4MemoryIF_M_AXI_ARVALID),
        .axi4MemoryIF_M_AXI_ARREADY (axi4MemoryIF_M_AXI_ARREADY),
        .axi4MemoryIF_M_AXI_RID (axi4MemoryIF_M_AXI_RID),
        .axi4MemoryIF_M_AXI_RDATA (axi4MemoryIF_M_AXI_RDATA),
        .axi4MemoryIF_M_AXI_RRESP (axi4MemoryIF_M_AXI_RRESP),
        .axi4MemoryIF_M_AXI_RLAST (axi4MemoryIF_M_AXI_RLAST),
        .axi4MemoryIF_M_AXI_RUSER (axi4MemoryIF_M_AXI_RUSER),
        .axi4MemoryIF_M_AXI_RVALID (axi4MemoryIF_M_AXI_RVALID),
        .axi4MemoryIF_M_AXI_RREADY (axi4MemoryIF_M_AXI_RREADY),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ACLK (axi4LitePlToPsControlRegisterIF_S_AXI_ACLK),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARESETN (axi4LitePlToPsControlRegisterIF_S_AXI_ARESETN),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARADDR (axi4LitePlToPsControlRegisterIF_S_AXI_ARADDR),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARPROT (axi4LitePlToPsControlRegisterIF_S_AXI_ARPROT),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARVALID (axi4LitePlToPsControlRegisterIF_S_AXI_ARVALID),
        .axi4LitePlToPsControlRegisterIF_S_AXI_ARREADY (axi4LitePlToPsControlRegisterIF_S_AXI_ARREADY),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RDATA (axi4LitePlToPsControlRegisterIF_S_AXI_RDATA),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RRESP (axi4LitePlToPsControlRegisterIF_S_AXI_RRESP),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RVALID (axi4LitePlToPsControlRegisterIF_S_AXI_RVALID),
        .axi4LitePlToPsControlRegisterIF_S_AXI_RREADY (axi4LitePlToPsControlRegisterIF_S_AXI_RREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ACLK (axi4LitePsToPlControlRegisterIF_S_AXI_ACLK),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARESETN (axi4LitePsToPlControlRegisterIF_S_AXI_ARESETN),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWADDR (axi4LitePsToPlControlRegisterIF_S_AXI_AWADDR),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWPROT (axi4LitePsToPlControlRegisterIF_S_AXI_AWPROT),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWVALID (axi4LitePsToPlControlRegisterIF_S_AXI_AWVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_AWREADY (axi4LitePsToPlControlRegisterIF_S_AXI_AWREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WDATA (axi4LitePsToPlControlRegisterIF_S_AXI_WDATA),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WSTRB (axi4LitePsToPlControlRegisterIF_S_AXI_WSTRB),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WVALID (axi4LitePsToPlControlRegisterIF_S_AXI_WVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_WREADY (axi4LitePsToPlControlRegisterIF_S_AXI_WREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_BRESP (axi4LitePsToPlControlRegisterIF_S_AXI_BRESP),
        .axi4LitePsToPlControlRegisterIF_S_AXI_BVALID (axi4LitePsToPlControlRegisterIF_S_AXI_BVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_BREADY (axi4LitePsToPlControlRegisterIF_S_AXI_BREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARADDR (axi4LitePsToPlControlRegisterIF_S_AXI_ARADDR),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARPROT (axi4LitePsToPlControlRegisterIF_S_AXI_ARPROT),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARVALID (axi4LitePsToPlControlRegisterIF_S_AXI_ARVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_ARREADY (axi4LitePsToPlControlRegisterIF_S_AXI_ARREADY),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RDATA (axi4LitePsToPlControlRegisterIF_S_AXI_RDATA),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RRESP (axi4LitePsToPlControlRegisterIF_S_AXI_RRESP),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RVALID (axi4LitePsToPlControlRegisterIF_S_AXI_RVALID),
        .axi4LitePsToPlControlRegisterIF_S_AXI_RREADY (axi4LitePsToPlControlRegisterIF_S_AXI_RREADY)
    );

endmodule : RSD
